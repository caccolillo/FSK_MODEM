library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity sinewave_generator is
    Port (
        clk               : in  std_logic;
        frequency_setting : in  std_logic_vector(7 downto 0); -- 8-bit frequency control
        sine_out          : out std_logic_vector(15 downto 0) -- 16-bit sine wave output
    );
end sinewave_generator;

architecture Behavioral of sinewave_generator is

    -- Constants
    constant LUT_SIZE : integer := 256;




  type sine_table_type is array(0 to 255) of unsigned(15 downto 0);

  signal sine_table : sine_table_type := (
      0 => to_unsigned(35446, 16),
      1 => to_unsigned(36182, 16),
      2 => to_unsigned(36918, 16),
      3 => to_unsigned(37652, 16),
      4 => to_unsigned(38385, 16),
      5 => to_unsigned(39118, 16),
      6 => to_unsigned(39847, 16),
      7 => to_unsigned(40574, 16),
      8 => to_unsigned(41298, 16),
      9 => to_unsigned(42019, 16),
     10 => to_unsigned(42735, 16),
     11 => to_unsigned(43447, 16),
     12 => to_unsigned(44154, 16),
     13 => to_unsigned(44855, 16),
     14 => to_unsigned(45551, 16),
     15 => to_unsigned(46241, 16),
     16 => to_unsigned(46924, 16),
     17 => to_unsigned(47602, 16),
     18 => to_unsigned(48271, 16),
     19 => to_unsigned(48933, 16),
     20 => to_unsigned(49586, 16),
     21 => to_unsigned(50232, 16),
     22 => to_unsigned(50868, 16),
     23 => to_unsigned(51494, 16),
     24 => to_unsigned(52111, 16),
     25 => to_unsigned(52718, 16),
     26 => to_unsigned(53314, 16),
     27 => to_unsigned(53899, 16),
     28 => to_unsigned(54473, 16),
     29 => to_unsigned(55035, 16),
     30 => to_unsigned(55586, 16),
     31 => to_unsigned(56123, 16),
     32 => to_unsigned(56658, 16),
     33 => to_unsigned(57178, 16),
     34 => to_unsigned(57687, 16),
     35 => to_unsigned(58182, 16),
     36 => to_unsigned(58663, 16),
     37 => to_unsigned(59130, 16),
     38 => to_unsigned(59583, 16),
     39 => to_unsigned(60012, 16),
     40 => to_unsigned(60427, 16),
     41 => to_unsigned(60826, 16),
     42 => to_unsigned(61209, 16),
     43 => to_unsigned(61577, 16),
     44 => to_unsigned(61929, 16),
     45 => to_unsigned(62265, 16),
     46 => to_unsigned(62583, 16),
     47 => to_unsigned(62887, 16),
     48 => to_unsigned(63172, 16),
     49 => to_unsigned(63440, 16),
     50 => to_unsigned(63691, 16),
     51 => to_unsigned(63925, 16),
     52 => to_unsigned(64141, 16),
     53 => to_unsigned(64338, 16),
     54 => to_unsigned(64519, 16),
     55 => to_unsigned(64690, 16),
     56 => to_unsigned(64852, 16),
     57 => to_unsigned(64997, 16),
     58 => to_unsigned(65122, 16),
     59 => to_unsigned(65229, 16),
     60 => to_unsigned(65327, 16),
     61 => to_unsigned(65406, 16),
     62 => to_unsigned(65466, 16),
     63 => to_unsigned(65508, 16),
     64 => to_unsigned(65531, 16),
     65 => to_unsigned(65535, 16),
     66 => to_unsigned(65520, 16),
     67 => to_unsigned(65486, 16),
     68 => to_unsigned(65434, 16),
     69 => to_unsigned(65363, 16),
     70 => to_unsigned(65273, 16),
     71 => to_unsigned(65165, 16),
     72 => to_unsigned(65038, 16),
     73 => to_unsigned(64892, 16),
     74 => to_unsigned(64728, 16),
     75 => to_unsigned(64546, 16),
     76 => to_unsigned(64346, 16),
     77 => to_unsigned(64127, 16),
     78 => to_unsigned(63890, 16),
     79 => to_unsigned(63634, 16),
     80 => to_unsigned(63361, 16),
     81 => to_unsigned(63069, 16),
     82 => to_unsigned(62759, 16),
     83 => to_unsigned(62432, 16),
     84 => to_unsigned(62087, 16),
     85 => to_unsigned(61725, 16),
     86 => to_unsigned(61345, 16),
     87 => to_unsigned(60948, 16),
     88 => to_unsigned(60535, 16),
     89 => to_unsigned(60103, 16),
     90 => to_unsigned(59656, 16),
     91 => to_unsigned(59193, 16),
     92 => to_unsigned(58712, 16),
     93 => to_unsigned(58216, 16),
     94 => to_unsigned(57703, 16),
     95 => to_unsigned(57176, 16),
     96 => to_unsigned(56632, 16),
     97 => to_unsigned(56073, 16),
     98 => to_unsigned(55500, 16),
     99 => to_unsigned(54912, 16),
    100 => to_unsigned(54308, 16),
    101 => to_unsigned(53690, 16),
    102 => to_unsigned(53059, 16),
    103 => to_unsigned(52413, 16),
    104 => to_unsigned(51753, 16),
    105 => to_unsigned(51079, 16),
    106 => to_unsigned(50393, 16),
    107 => to_unsigned(49693, 16),
    108 => to_unsigned(48980, 16),
    109 => to_unsigned(48255, 16),
    110 => to_unsigned(47517, 16),
    111 => to_unsigned(46768, 16),
    112 => to_unsigned(46007, 16),
    113 => to_unsigned(45235, 16),
    114 => to_unsigned(44461, 16),
    115 => to_unsigned(43675, 16),
    116 => to_unsigned(42879, 16),
    117 => to_unsigned(42082, 16),
    118 => to_unsigned(41284, 16),
    119 => to_unsigned(40485, 16),
    120 => to_unsigned(39684, 16),
    121 => to_unsigned(38884, 16),
    122 => to_unsigned(38084, 16),
    123 => to_unsigned(37284, 16),
    124 => to_unsigned(36484, 16),
    125 => to_unsigned(35685, 16),
    126 => to_unsigned(34885, 16),
    127 => to_unsigned(34086, 16),
    128 => to_unsigned(33287, 16),
    129 => to_unsigned(32489, 16),
    130 => to_unsigned(31690, 16),
    131 => to_unsigned(30894, 16),
    132 => to_unsigned(30099, 16),
    133 => to_unsigned(29307, 16),
    134 => to_unsigned(28516, 16),
    135 => to_unsigned(27728, 16),
    136 => to_unsigned(26944, 16),
    137 => to_unsigned(26162, 16),
    138 => to_unsigned(25384, 16),
    139 => to_unsigned(24610, 16),
    140 => to_unsigned(23841, 16),
    141 => to_unsigned(23077, 16),
    142 => to_unsigned(22318, 16),
    143 => to_unsigned(21564, 16),
    144 => to_unsigned(20818, 16),
    145 => to_unsigned(20078, 16),
    146 => to_unsigned(19346, 16),
    147 => to_unsigned(18621, 16),
    148 => to_unsigned(17905, 16),
    149 => to_unsigned(17197, 16),
    150 => to_unsigned(16499, 16),
    151 => to_unsigned(15810, 16),
    152 => to_unsigned(15130, 16),
    153 => to_unsigned(14462, 16),
    154 => to_unsigned(13805, 16),
    155 => to_unsigned(13157, 16),
    156 => to_unsigned(12523, 16),
    157 => to_unsigned(11899, 16),
    158 => to_unsigned(11289, 16),
    159 => to_unsigned(10690, 16),
    160 => to_unsigned(10105, 16),
    161 => to_unsigned(9533, 16),
    162 => to_unsigned(8975, 16),
    163 => to_unsigned(8430, 16),
    164 => to_unsigned(7900, 16),
    165 => to_unsigned(7384, 16),
    166 => to_unsigned(6884, 16),
    167 => to_unsigned(6398, 16),
    168 => to_unsigned(5929, 16),
    169 => to_unsigned(5475, 16),
    170 => to_unsigned(5037, 16),
    171 => to_unsigned(4616, 16),
    172 => to_unsigned(4211, 16),
    173 => to_unsigned(3824, 16),
    174 => to_unsigned(3453, 16),
    175 => to_unsigned(3101, 16),
    176 => to_unsigned(2766, 16),
    177 => to_unsigned(2448, 16),
    178 => to_unsigned(2150, 16),
    179 => to_unsigned(1869, 16),
    180 => to_unsigned(1608, 16),
    181 => to_unsigned(1366, 16),
    182 => to_unsigned(1143, 16),
    183 => to_unsigned(938, 16),
    184 => to_unsigned(754, 16),
    185 => to_unsigned(590, 16),
    186 => to_unsigned(446, 16),
    187 => to_unsigned(321, 16),
    188 => to_unsigned(217, 16),
    189 => to_unsigned(133, 16),
    190 => to_unsigned(70, 16),
    191 => to_unsigned(26, 16),
    192 => to_unsigned(3, 16),
    193 => to_unsigned(0, 16),
    194 => to_unsigned(18, 16),
    195 => to_unsigned(57, 16),
    196 => to_unsigned(116, 16),
    197 => to_unsigned(196, 16),
    198 => to_unsigned(297, 16),
    199 => to_unsigned(418, 16),
    200 => to_unsigned(560, 16),
    201 => to_unsigned(723, 16),
    202 => to_unsigned(907, 16),
    203 => to_unsigned(1112, 16),
    204 => to_unsigned(1338, 16),
    205 => to_unsigned(1584, 16),
    206 => to_unsigned(1851, 16),
    207 => to_unsigned(2139, 16),
    208 => to_unsigned(2448, 16),
    209 => to_unsigned(2778, 16),
    210 => to_unsigned(3128, 16),
    211 => to_unsigned(3499, 16),
    212 => to_unsigned(3891, 16),
    213 => to_unsigned(4303, 16),
    214 => to_unsigned(4735, 16),
    215 => to_unsigned(5188, 16),
    216 => to_unsigned(5661, 16),
    217 => to_unsigned(6155, 16),
    218 => to_unsigned(6668, 16),
    219 => to_unsigned(7201, 16),
    220 => to_unsigned(7754, 16),
    221 => to_unsigned(8327, 16),
    222 => to_unsigned(8920, 16),
    223 => to_unsigned(9531, 16),
    224 => to_unsigned(10163, 16),
    225 => to_unsigned(10813, 16),
    226 => to_unsigned(11482, 16),
    227 => to_unsigned(12170, 16),
    228 => to_unsigned(12878, 16),
    229 => to_unsigned(13604, 16),
    230 => to_unsigned(14349, 16),
    231 => to_unsigned(15113, 16),
    232 => to_unsigned(15895, 16),
    233 => to_unsigned(16695, 16),
    234 => to_unsigned(17513, 16),
    235 => to_unsigned(18349, 16),
    236 => to_unsigned(19203, 16),
    237 => to_unsigned(20075, 16),
    238 => to_unsigned(20964, 16),
    239 => to_unsigned(21870, 16),
    240 => to_unsigned(22794, 16),
    241 => to_unsigned(23734, 16),
    242 => to_unsigned(24692, 16),
    243 => to_unsigned(25666, 16),
    244 => to_unsigned(26658, 16),
    245 => to_unsigned(27666, 16),
    246 => to_unsigned(28689, 16),
    247 => to_unsigned(29730, 16),
    248 => to_unsigned(30787, 16),
    249 => to_unsigned(31860, 16),
    250 => to_unsigned(32949, 16),
    251 => to_unsigned(34054, 16),
    252 => to_unsigned(35174, 16),
    253 => to_unsigned(36308, 16),
    254 => to_unsigned(37459, 16),
    255 => to_unsigned(38615, 16)
  );



    -- Internal signals
    signal phase_accumulator : unsigned(15 downto 0) := (others => '0');
    signal phase_increment   : unsigned(15 downto 0);

begin

    -- Calculate phase increment from frequency setting
    process(frequency_setting)
    begin
        -- Map 8-bit frequency setting to 16-bit phase increment
        -- Simple linear mapping: frequency_setting * constant
        phase_increment <= resize(unsigned(frequency_setting) * 4, 16);  -- Scale factor is arbitrary
    end process;

    -- Phase accumulator and LUT access
    process(clk)
    begin
        if rising_edge(clk) then
            phase_accumulator <= phase_accumulator + phase_increment;
        end if;
    end process;

    -- Output sine wave sample from LUT
    sine_out <= std_logic_vector(sine_table(to_integer(phase_accumulator(15 downto 8))));

end Behavioral;

